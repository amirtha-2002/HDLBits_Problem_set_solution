module top_module( 
    input a, 
    input b, 
    output out );
    and g1(out,a,b);

endmodule
