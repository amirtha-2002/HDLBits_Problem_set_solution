module top_module( 
    input a, 
    input b, 
    output out );
    nor g1(out,a,b);

endmodule
